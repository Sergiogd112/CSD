--------------------------------------------------------------------------------
-- An example of a 4-bit full adder (Adder_4bit) using a hierarchical structure
-- This VHDL file is a translation of the following schematic:
-- https://digsys.upc.edu/csd/P03/P3_T/Plan_PC_Adder_4bit_ripple_carry.pdf
---------------------------------------------------
-- This example file can be used as a seed to copy and adapt any other 
-- hiearchical design based on components and signals 
---------------------------------------------------
-- Exercise P3  - CSD - Arithmetic circuits
-- http://digsys.upc.edu
--------------------------------------------------------------------------------

LIBRARY ieee;
USE  IEEE.STD_LOGIC_1164.all;

ENTITY Adder_4bit IS

	PORT (
		A,B	: IN 	STD_LOGIC_VECTOR(3 DOWNTO 0); 				
		Cin	: IN 	STD_LOGIC;    
		S	: OUT 	STD_LOGIC_VECTOR (3 DOWNTO 0);
		Cout	: OUT  	STD_LOGIC;
		Z	: OUT 	STD_LOGIC		-- Z = 0 when S(3..0) and  C4 = 0;
	  );

END Adder_4bit;


ARCHITECTURE hierarchical_structure OF Adder_4bit IS

	
-- The elemental component to be used:
 
	COMPONENT Adder_1bit IS  

		PORT (
			Ai,Bi, Ci	: IN STD_LOGIC;				
			So, Co		: OUT STD_LOGIC
		  );

	END COMPONENT;

-- Signals

	SIGNAL	C1, C2, C3, C4 	: STD_LOGIC;	-- The wires to connect 1-bit modules together 
	SIGNAL	Y	 	: STD_LOGIC_VECTOR (3 DOWNTO 0);

BEGIN

-- Instantiation of up to 4 basic 1-bit adders:

	Chip0	: Adder_1bit
		PORT MAP (
	-- from component name 	=> to signal or port name
			Ai		=> A(0),
			Bi 		=> B(0),
			Ci 		=> Cin,
			So	 	=> Y(0), 
			Co	 	=> C1 					  
		);

	Chip1	: Adder_1bit
		PORT MAP (
				-- from component name 	=> to signal or port name
			Ai		=> A(1),
			Bi 		=> B(1),
			Ci 		=> C1,
			So	 	=> Y(1), 
			Co	 	=> C2 					  
		);

	Chip2	: Adder_1bit
		PORT MAP (
-- from component name 	=> to signal or port name
					Ai		=> A(2),
					Bi 		=> B(2),
					Ci 		=> C2,
					So	 	=> Y(2), 
					Co	 	=> C3 					  
		);

	Chip3	: Adder_1bit
		PORT MAP (
-- from component name 	=> to signal or port name
			Ai			=> A(3),
			Bi 			=> B(3),
			Ci 			=> C3,
			So	 		=> Y(3), 
			Co	 		=> C4 					  
		);

-- Other circuits and equations:

S <= Y;

Z <= NOT (Y(3) OR Y(2) OR Y(1) OR Y(0) OR C4 );

Cout <= C4;

			 		   	 		 		   	   
END hierarchical_structure;
